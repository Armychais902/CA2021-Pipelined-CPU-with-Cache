module EX_MEM
(
    clk_i,
	start_i,
	MemStall_i,
    RegWrite_i,
    MemtoReg_i,
    MemRead_i,
    MemWrite_i,
    ALUResult_i,
    RS2data_i,
	RDaddr_i,
	RegWrite_o,
	MemtoReg_o,
	MemRead_o,
	MemWrite_o,
	ALUResult_o,
	RS2data_o,
	RDaddr_o
);

input           clk_i;
input			start_i;
input 			MemStall_i;
input           RegWrite_i, MemtoReg_i, MemRead_i, MemWrite_i;
input [4:0]     RDaddr_i;
input [31:0]    ALUResult_i, RS2data_i;
output reg      RegWrite_o, MemtoReg_o, MemRead_o, MemWrite_o;
output	[4:0]   RDaddr_o;
reg		[4:0]   RDaddr_o;
output 	[31:0]  ALUResult_o, RS2data_o;
reg		[31:0]  ALUResult_o, RS2data_o;

always @(posedge clk_i or negedge start_i) begin
	if (!start_i)	begin
		RegWrite_o <= 1'b0;
		MemtoReg_o <= 1'b0;
		MemRead_o <= 1'b0;
		MemWrite_o <= 1'b0;
		ALUResult_o <= 32'b0;
		RS2data_o <= 32'b0;
		RDaddr_o <= 5'b0;
	end
	else if (!MemStall_i)	begin
		RegWrite_o <= RegWrite_i;
		MemtoReg_o <= MemtoReg_i;
		MemRead_o <= MemRead_i;
		MemWrite_o <= MemWrite_i;
		ALUResult_o <= ALUResult_i;
		RS2data_o <= RS2data_i;
		RDaddr_o <= RDaddr_i;
	end
end

endmodule